module obstacle_control (
    input clk,
    input speed,
    input en1,
    output reg [9:0] hCount1,
    output reg [9:0] hCount2,
    output reg [9:0] hCount3,
);

//local variable
reg [2:0] num_obs;

always @(posedge clk ) begin

    
end
    
endmodule